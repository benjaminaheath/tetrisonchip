module test_piecegenerator;


endmodule
