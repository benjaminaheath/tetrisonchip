`include "include/part.sv"
module chip(

);

board_mem prev_state(.*);
board_mem curr_state(.*);

endmodule