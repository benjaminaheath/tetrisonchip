module chip(

);

board prev_state(.*);
board curr_state(.*);

endmodule