typedef struct {
    logic filled;
    logic active;
} tile;